module tb();
reg [15:0]A;
reg [15:0]B;
reg cin;
wire [15:0]sum;
wire cout;

Select_Carry_Adder sC (A,B,cin,cout,sum); 
initial begin
$monitor("Time=%g",$time,"A=%b,B=%b,Cin=%b : Sum= %b,Cout=%b",A,B,cin,sum,cout);
 A= 16'b0000000000011111; B=16'b000000000001100; cin=1'b0;
#10  A= 16'b1100011000011111; B=16'b000000110001100; cin=1'b1;
#10 A= 16'b1111111111111111; B=16'b000000000000000; cin=1'b1;
#10 A= 16'b1001001001001001; B=16'b1001001001001001; cin=1'b1;
end
endmodule


//////////////////
output
Time=0A=0000000000011111,B=0000000000001100,Cin=0 : Sum= 0000000000101011,Cout=0
Time=10A=1100011000011111,B=0000000110001100,Cin=1 : Sum= 1100011110101100,Cout=0
Time=20A=1111111111111111,B=0000000000000000,Cin=1 : Sum= 0000000000000000,Cout=1
Time=30A=1001001001001001,B=1001001001001001,Cin=1 : Sum= 0010010010010011,Cout=1
